`timescale 1ns / 1ps

module pulse_controller (
    input clk,
    input sw_input,
    input clear,
    output logic clk_pulse
);

  logic [2:0] state, nextstate;
  logic [27:0] CNT;
  wire cnt_zero;

  always @(posedge clk, posedge clear)
    if (clear) state <= 3'b000;
    else state <= nextstate;

  always @(sw_input, state, cnt_zero)
    case (state)
      3'b000: begin
        if (sw_input) nextstate = 3'b001;
        else nextstate = 3'b000;
        clk_pulse = 0;
      end
      3'b001: begin
        nextstate = 3'b010;
        clk_pulse = 1;
      end
      3'b010: begin
        if (cnt_zero) nextstate = 3'b011;
        else nextstate = 3'b010;
        clk_pulse = 1;
      end
      3'b011: begin
        if (sw_input) nextstate = 3'b011;
        else nextstate = 3'b100;
        clk_pulse = 0;
      end
      3'b100: begin
        if (cnt_zero) nextstate = 3'b000;
        else nextstate = 3'b100;
        clk_pulse = 0;
      end
      default: begin
        nextstate = 3'b000;
        clk_pulse = 0;
      end
    endcase

  always @(posedge clk)
    unique case (state)
      3'b001: CNT <= 100000000;
      3'b010: CNT <= CNT - 1;
      3'b011: CNT <= 100000000;
      3'b100: CNT <= CNT - 1;
    endcase

  // reduction operator |CNT gives the OR of all bits in the CNT register
  assign cnt_zero = ~|CNT;

endmodule
