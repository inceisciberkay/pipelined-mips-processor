`timescale 1ns / 1ps

module mips (
    input logic clk,
    input logic reset,
    output logic [31:0] pc,
    output logic [31:0] pcn,
    input logic [31:0] instrF,
    output logic MemWriteM,
    output logic [31:0] ALUOutM,
    output logic [31:0] resultW,
    output logic [31:0] instrOut,
    input logic [31:0] ReadDataM,
    output logic [31:0] WriteDataM,
    output logic ZeroM,
    output logic BranchM,
    output logic ZeroE,
    output logic RegWriteE,
    output logic MemtoRegE,
    output logic MemWriteE,
    output logic [31:0] SrcAE,
    output logic [31:0] SrcBE,
    output logic [31:0] ALUOutE,
    output logic [31:0] WriteDataE,
    output logic BranchE,
    output logic [4:0] WriteRegE,
    output logic [31:0] PCBranchE,
    output logic [31:0] instrD,
    output logic [31:0] instrE,
    output logic [31:0] instrM,
    output logic [31:0] instrW,
    output logic [1:0] ForwardAE,
    output logic [1:0] ForwardBE,
    output logic [31:0] RD1E,
    output logic [31:0] RD2E,
    output logic [31:0] RD1,
    output logic [31:0] RD2,
    output logic ALUSrcE,
    output logic [31:0] SignImmE,
    output logic [31:0] PCBranchM
);

  logic MemWriteD, MemToRegD, pcsrc, zero, ALUSrcD, RegDstD, RegWriteD, BranchD;
  logic [2:0] ALUControlD;
  assign instrOut = instrF;
  logic Jump;

  controller c (
      .op(instrD[31:26]),
      .funct(instrD[5:0]),
      .memtoreg(MemToRegD),
      .memwrite(MemWriteD),
      .alusrc(ALUSrcD),
      .regdst(RegDstD),
      .regwrite(RegWriteD),
      .jump(Jump),
      .alucontrol(ALUControlD),
      .branch(BranchD)
  );

  datapath dp (
      .clk(clk),
      .reset(reset),
      .RegWriteD(RegWriteD),
      .MemtoRegD(MemToRegD),
      .MemWriteD(MemWriteD),
      .ALUSrcD(ALUSrcD),
      .RegDstD(RegDstD),
      .ALUControlD(ALUControlD),
      .BranchD(BranchD),
      .rsD(instrD[25:21]),
      .rtD(instrD[20:16]),
      .rdD(instrD[15:11]),
      .immD(instrD[15:0]),
      .instrF(instrF),
      .PCF(pc),
      .PCN(pcn),
      .instrD(instrD),
      .MemWriteM(MemWriteM),
      .ALUOutM(ALUOutM),
      .ReadDataM(ReadDataM),
      .Jump(Jump),
      .WriteDataM(WriteDataM),
      .ZeroM(ZeroM),
      .BranchM(BranchM),
      .ZeroE(ZeroE),
      .RegWriteE(RegWriteE),
      .MemtoRegE(MemtoRegE),
      .MemWriteE(MemWriteE),
      .SrcAE(SrcAE),
      .SrcBE(SrcBE),
      .ALUOutE(ALUOutE),
      .WriteDataE(WriteDataE),
      .BranchE(BranchE),
      .WriteRegE(WriteRegE),
      .PCBranchE(PCBranchE),
      .instrE(instrE),
      .instrM(instrM),
      .instrW(instrW),
      .ForwardAE(ForwardAE),
      .ForwardBE(ForwardBE),
      .RD1E(RD1E),
      .RD2E(RD2E),
      .RD1(RD1),
      .RD2(RD2),
      .ALUSrcE(ALUSrcE),
      .SignImmE(SignImmE),
      .PCBranchM(PCBranchM)
  );

endmodule
