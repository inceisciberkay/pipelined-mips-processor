`timescale 1ns / 1ps

module PipeWtoF (
    input logic [31:0] PC,
    input logic EN,
    input logic clk,
    input logic reset,  // StallF will be connected as this EN
    output logic [31:0] PCF
);

  always_ff @(posedge clk, posedge reset)
    if (reset) PCF <= 0;
    else if (EN) PCF <= PC;

endmodule
